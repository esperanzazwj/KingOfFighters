`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:16:11 01/08/2016 
// Design Name: 
// Module Name:    bg_rom_g 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module bg_rom_g(input wire clk, input wire[6:0] addr, output reg[159:0] bitmap);
	reg [6:0] addr_reg;
	always @(posedge clk)
		addr_reg<=addr;
	always @(*)
	begin
		case (addr_reg)
7'd000:bitmap<=160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd001:bitmap<=160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd002:bitmap<=160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd003:bitmap<=160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd004:bitmap<=160'b1111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd005:bitmap<=160'b1111111111111111111111111111111111111111111111111111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd006:bitmap<=160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd007:bitmap<=160'b1111111111111110111111111111111111111111111111111111110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd008:bitmap<=160'b1111111111111110011111111111111111111111111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd009:bitmap<=160'b1111111111111100101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd010:bitmap<=160'b1111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd011:bitmap<=160'b1111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd012:bitmap<=160'b1111111111110011111111011111111111111111111111111111011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd013:bitmap<=160'b1111111111100001011111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd014:bitmap<=160'b1111111111101011111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd015:bitmap<=160'b1111111111111111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111000100;
7'd016:bitmap<=160'b1111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110000011111111;
7'd017:bitmap<=160'b1111111111111111111101111111110111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd018:bitmap<=160'b1111111111111111111111101111111001111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd019:bitmap<=160'b1111111111111111111111111111111110111111110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd020:bitmap<=160'b1111111111111111111111111111111111111111110000110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd021:bitmap<=160'b1111111111111111111111111111111111110111110100110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd022:bitmap<=160'b1111111111111111111111111111110111111101111110101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd023:bitmap<=160'b1111111111111111111111111111111011111110100001101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd024:bitmap<=160'b1111111111111111111111111111111110111111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd025:bitmap<=160'b1111111111111111111111111111111111100111110010011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd026:bitmap<=160'b1111111111111111111111111111111111111001101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd027:bitmap<=160'b1111111111111111111111111111111111111110001111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd028:bitmap<=160'b1111111111111111111111111111111111111111000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd029:bitmap<=160'b1111111111111111111111111111111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd030:bitmap<=160'b1111111111111111111111111111111111111100010000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd031:bitmap<=160'b1111111111111111111111111111111111111110010000000101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd032:bitmap<=160'b1111111111111111111111111111111111111110100100000111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111;
7'd033:bitmap<=160'b1111111111111111111111111111111111111110011000000111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd034:bitmap<=160'b1111111111111111111111111111111111111110011100001111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111;
7'd035:bitmap<=160'b1111111111111111111111111111111111111110111000001111111111011111111111111111111111111111111111111111111111111111111111111111111101111111111111111110101110111111;
7'd036:bitmap<=160'b1111111111111111111111111111111111111111111000011111011111110111111111111111111111111111111111111111111111111111111111111111110111111111111111111110110011100111;
7'd037:bitmap<=160'b1111111111111111111111111111111111111111111100011111111111111101111111111111111111111111111111111111111111111111111111111111011111111111111111111111000011101101;
7'd038:bitmap<=160'b1111111111111111111111111111111111111111110000011111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111100111110110001010;
7'd039:bitmap<=160'b1111111111111111111111111111111111111111111100011111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111110110111100000000;
7'd040:bitmap<=160'b1111111111111111111111111111111111110111101110011111111111111111111101111111111111111111111111111111111111111111111111111101111111111111111111101110110000001000;
7'd041:bitmap<=160'b1111111111111111111111111111111111111111110010111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111101110000101000100;
7'd042:bitmap<=160'b1111111111111111111111111111111111101111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000010000;
7'd043:bitmap<=160'b1111111111111111111111111111111111001111000011111111111111111111001111101101111111111111111111111111111111111111111111111111111111111111111111111110000000011000;
7'd044:bitmap<=160'b1111111111111111111111111110111111011111000011111111111111111111111111111110111111111111111111111111111111111111111111100111111111111111111111111111100000000000;
7'd045:bitmap<=160'b1111111111111111111111111111111111111110000111111111111111111111111111011011111111111111111111111111111111111111111111100111111111111111111111111111110001010000;
7'd046:bitmap<=160'b1111111111111111111111111111111110111110000111111111111111111111111110010001111111111111111111111111111111111111111111111111111111111111111111111111111000010000;
7'd047:bitmap<=160'b1111111111111111111111111111111111111110000111111111111111111111111111000101111111111111111111111111111111111111111100111111111111111111111111111111111111000000;
7'd048:bitmap<=160'b1111111111111111111111100111111101111101001111111111111111111111111111100011111111111111111111111111111111111111101111111111111111111111111111111111111111110000;
7'd049:bitmap<=160'b1111111111111111111111110001111011111101000111111111111111111111111111000001111111111111111111111111111111111111000011111111111111111111111111111111111111111110;
7'd050:bitmap<=160'b1111111111111111111111111011111111111111001111111111111111111111111111101010111111111111111110011111111111111111111101111111111111111111111111111111111111111111;
7'd051:bitmap<=160'b1111111111111111101111111011110111111010001111111111111111111111111111110011111111111111111100011111111111111111111111111111111111110111111111111111111111111111;
7'd052:bitmap<=160'b1111111111111111111111000111110111111010001111111111111111111111111111100011011111111111101100011111111111111111011101111111111111111111111111111111111111111111;
7'd053:bitmap<=160'b1111111111111110111111110111101111111110001111111111111111111111111110100001011011111111100111111111111111111111001110111111111111111111111111111111111111111111;
7'd054:bitmap<=160'b1111111111111111111111111011011111010100001111111111111111111111111111001000011111111111011111111011111111111111100001110111111111111111111111111111111111111111;
7'd055:bitmap<=160'b1110100010101111100111100101101111110100010000111111111111111110001111011111000111110110001111111101111111111101111111111111111111111111111111111111111111111111;
7'd056:bitmap<=160'b1111111000011111101111011101111111110000000000110111111111111110000011100100001100110011001111111000111111110111111111111111111111111111111111111111111111111111;
7'd057:bitmap<=160'b1111110101011111101110000011110111110000000000000011111111111101000011000000001010110111011111111110111110111111111111101111111111111111111111111111111111111110;
7'd058:bitmap<=160'b1101010100001111110110000111011111111110000000000111111111100000000111000010000000000100011011111111111111011111111111111111111111111111111111111111111111111100;
7'd059:bitmap<=160'b1101110010011111111110010010111111110100001110000111111111110000001000000011000001000000000001111111111101011110111111111111111111111111111111111111111111110000;
7'd060:bitmap<=160'b1101011010111111101100111111110111111000000001001111110111101000000000000001100000000000000001111111111100011000111111111111111111111111111111111111111111110000;
7'd061:bitmap<=160'b1000110111111101111111110110010110110000000100000111111111101100000000010011110000000000000000111111110000111110001111111111111111111111111111111111111111100000;
7'd062:bitmap<=160'b1100001111111101000010000000000001110100111100001111111111111100000000010011100000000000000000111111100000110010011111111111110111111111111111111111111111000011;
7'd063:bitmap<=160'b0000001111110000001100011000000000001101111111001111111111111100000000010011100000000000000000111101100000111010011111111111111111110101010011111111111110001111;
7'd064:bitmap<=160'b0000000011000000000011101100000000000001111111110001111110000000000000000011100000000001000000001110100000111010011111100010110111110100000001001111111011111111;
7'd065:bitmap<=160'b1100001000111000001111111000000000000000011111000111111110100000000000010000000000000000000000011000000000010000111101101000110101100000000000011111110111111111;
7'd066:bitmap<=160'b1011000000000000011111111000010110000001100110111100000000000000000000111011000000000000000000011011110000011001111101100001100011100000000000011111111111111111;
7'd067:bitmap<=160'b1100000010101010110111110000000000000111111111111011111100000000000011001110000000000011000000011111110000011111111101100000100000000000000000011111101000001111;
7'd068:bitmap<=160'b1100000001100101111111110000000000000000000000000011111101101000000000000000000000000111000000001111111111111111111011000000101000000000000000001101000000001000;
7'd069:bitmap<=160'b0101010100010111111111000000000000000000000000000000000110100011100000001100000110001111000110000101111111111111111001000000100000000000000000000000000000000000;
7'd070:bitmap<=160'b1111010010111111111110000000001111110000000000000011111111111111010000001000001111001111100111000011001111111111111000000000100100000000000000000000000000000000;
7'd071:bitmap<=160'b1000000011111111111100000011111111111111000000000001111111011101010000000000011100000001100110001001111011111110011000000000100000000000000000000000011000000000;
7'd072:bitmap<=160'b0101011111111111111100001111111111111111110000000001111111111110000000000011111100000000100010000011110011111000011001100000110100000000000000000000011000000000;
7'd073:bitmap<=160'b1001111111111111100000001010011111111111111000001011111111110000000000001011111110000011100010110000110111111000011111100000111000000000000000000000000000000000;
7'd074:bitmap<=160'b0100111011000010000000000001110111101111011110000011111111111001000000000111111111000011100000001000110111111000111111100000111000000000000000000011000000000000;
7'd075:bitmap<=160'b0000000000000000000000101001001110111001111000101111110000111110000000000001111111100000000001010101100111111000011010100000110000000000000000000111111000000000;
7'd076:bitmap<=160'b0000000000000000000000010000101011111111100000000010000000000000000101000000001000000011000000001100100000001011111101101110110011000000000100000111111000000000;
7'd077:bitmap<=160'b0000000000000000000000100101101111000010000000000000001110000000000000000000000000000001110001001111100000011111111111111111111010000000001110111111111100000000;
7'd078:bitmap<=160'b0000000000000000000000000000001010100000000000000000001010000000000000000000000000000011010000001011100000001111111100111111111110000000000011111111111100000001;
7'd079:bitmap<=160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000011101111000001111111011110000111111111000101011111111110000000000;
7'd080:bitmap<=160'b0000000000000000000000000000000000000000000000000000011110110000001000000000000000000010010000011111101000001110110111100000000111111111111111111111110000000000;
7'd081:bitmap<=160'b0000000000000000000000000000000000000000000000000000001110000000000000000000000000001111111000011111111111110111000011100000101011111111111111111011110000000000;
7'd082:bitmap<=160'b0000000000000000000000000000000000000000000000000000001110000000001101101000000000111111110000011111101111111111111111111111110111111111111111111101111110000000;
7'd083:bitmap<=160'b1111100000000000000000000000000000000000000000000000011110100000000000000000000001111111100001111111111111111111111111111111111111111111111111111100011100000000;
7'd084:bitmap<=160'b1111100000000001000000000000000000000000000000000100001110001001000000000001101011111111100111111111101111111111111111111111111111111111111111111110001100000000;
7'd085:bitmap<=160'b1111111100000000110000000000000000000000000000000100011111111010000001000011111111110011000111111111101111111111111111111111111111111111111111111111000000000000;
7'd086:bitmap<=160'b1111111100000001100000000000000000000000000000001101111111111111100000001111110010100101000111111111100001111111111111111111111111111111111111111111000000000000;
7'd087:bitmap<=160'b1110111110000001110000000000000000000000000000001001011111111100000000111111100001000001000111111011100000111111111111111111111111111111111111111111000000000000;
7'd088:bitmap<=160'b1000111100000001100000000000000000000000000010001111111111111000000111111111100000000010001100000001000001111111111111111111111111111100111111111111000000000000;
7'd089:bitmap<=160'b0100111000000001000000000000000000000000000010001111111111111011111111111111100000000010001000000001000011111111111111110111111111111100111111111000000000000000;
7'd090:bitmap<=160'b0000011000000001100000000000000000000000000000011111111111111111100010111111000000000010000011110000000000010111111111100111111111110001111111111100000000000000;
7'd091:bitmap<=160'b0010000000000000100000000000000000000000000100111111111111111111111111111111000000000010000001110000000000000011111100010111111111110000011111101000000000000000;
7'd092:bitmap<=160'b0000100000000000100000000000000000000000101111111111111111111111111101111111010000000000000000100000000000000110000000001000111110000000001111111100000000000000;
7'd093:bitmap<=160'b0101000000000000100000000000000010011111111111111111111111111111111111111111111000000110110000100010000000001100000101111111101111000000000011111100000000000000;
7'd094:bitmap<=160'b1010000000000000100000000000000011000000011110001111111111111111111111111111111000000000110010011101000000000001001011111011111100110000000001001110111000000000;
7'd095:bitmap<=160'b1000000000000000000000000000000011000000000000001011111111111111111111111111111110100000011110001110000000000000110111110111110001110000000000011100111100000000;
7'd096:bitmap<=160'b0110000000000000000000000000000011000000000000001111111111111111111111111111011110000000001111000110000100000000000000101001000100110000000000011001111111000000;
7'd097:bitmap<=160'b1000000000000000100000000000000011000000000000001111111111111111111111111110001100000000001111111101000100000000000101000011000000000000000000010000011111101100;
7'd098:bitmap<=160'b0000000000000000100000000000000011000000000000001111111111111111111111111000000000000000000101111001100000000000100000111101110000111000000100000000010111110000;
7'd099:bitmap<=160'b0000000000000000100000000000000011000000000000001111111111111111111111110000000110000000001111111010100000000000010000001001101010001110000000000000000111111000;
7'd100:bitmap<=160'b0000000000000000100101000000000011000000000000000101111111111111111111111111111100000000001101111110000000000000100001111111111111110110100000000011000001111100;
7'd101:bitmap<=160'b0000000000000000000010100000000011000000000000000001111111111111111111111111111100000000000001100000000000000000001100111111111001111111111111001111111000011110;
7'd102:bitmap<=160'b1000000000000000011111110000000001000000000000000001111111111111111111111111111100000000000000000000000000000000111111111111111111111111011110111111111111111111;
7'd103:bitmap<=160'b0100000000000000011111100000000000000000000000010001111111111111111111111111111100111110000100000111000000110011111111111111111111111111111111111111111111111111;
7'd104:bitmap<=160'b1000000000000000001101100100000000001000000000000000111111111111111111111111111111111111111111111111110001111111111111111111111111111111111111111111111111111111;
7'd105:bitmap<=160'b0000000000000000000011010100000000000000000000001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd106:bitmap<=160'b0000000000000000000100000100000000000000000000111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd107:bitmap<=160'b0001000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd108:bitmap<=160'b0000111100000000000000011000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd109:bitmap<=160'b0001000000000000000000000100000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd110:bitmap<=160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd111:bitmap<=160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd112:bitmap<=160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd113:bitmap<=160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd114:bitmap<=160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd115:bitmap<=160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd116:bitmap<=160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd117:bitmap<=160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd118:bitmap<=160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd119:bitmap<=160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		
		endcase
	end
endmodule

`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:16:27 01/08/2016 
// Design Name: 
// Module Name:    bg_rom_b 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module bg_rom_b(input wire clk, input wire[6:0] addr, output reg[159:0] bitmap);
	reg [6:0] addr_reg;
	always @(posedge clk)
		addr_reg<=addr;
	always @(*)
	begin
		case (addr_reg)
7'd000:bitmap<=160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd001:bitmap<=160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd002:bitmap<=160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd003:bitmap<=160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd004:bitmap<=160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd005:bitmap<=160'b1111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd006:bitmap<=160'b1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd007:bitmap<=160'b1111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd008:bitmap<=160'b1111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd009:bitmap<=160'b1111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd010:bitmap<=160'b1111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd011:bitmap<=160'b1111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd012:bitmap<=160'b1111111111110011111111011111111111111111111111111111011110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd013:bitmap<=160'b1111111111100011111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000;
7'd014:bitmap<=160'b1111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111110100000000;
7'd015:bitmap<=160'b1111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000100;
7'd016:bitmap<=160'b1111111111111111111111111111011111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100110000000010111;
7'd017:bitmap<=160'b1111111111111111111101111111110111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd018:bitmap<=160'b1111111111111111111111111111111011111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd019:bitmap<=160'b1111111111111111111111111111111110111111110000011111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd020:bitmap<=160'b1111111111111111111111111111111111111111110000110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd021:bitmap<=160'b1111111111111111111111111111111111111111110000110111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd022:bitmap<=160'b1111111111111111111111111111110111111101110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd023:bitmap<=160'b1111111111111111111111111111111011111110110000101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd024:bitmap<=160'b1111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd025:bitmap<=160'b1111111111111111111111111111111111110111110110011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd026:bitmap<=160'b1111111111111111111111111111111111111101101111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd027:bitmap<=160'b1111111111111111111111111111111111111110001111011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd028:bitmap<=160'b1111111111111111111111111111111111111110000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd029:bitmap<=160'b1111111111111111111111111111111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd030:bitmap<=160'b1111111111111111111111111111111111111100010000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd031:bitmap<=160'b1111111111111111111111111111111111111110000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010111111111;
7'd032:bitmap<=160'b1111111111111111111111111111111111111110000000000011011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001111111;
7'd033:bitmap<=160'b1111111111111111111111111111111111111110011000000111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001000111111;
7'd034:bitmap<=160'b1111111111111111111111111111111111111110011100001011111101111111111111111111111111111111111111111111111111111111111111111111111000000111111111111100000000110101;
7'd035:bitmap<=160'b1111111111111111111111111111111111111110111000001111111111011111111111111111111111111111111111111111111111111111111111111111110000111111111111111100000000000001;
7'd036:bitmap<=160'b1111111111111111111111111111111111111111111000011111111111100111111111111111111111111111111111111111111111111111111111111111000111111111111111110000000000000000;
7'd037:bitmap<=160'b1111111111111111111111111111111111111111111001011111111111111101111111111111111111111111111111111111111111111111111111111110011111111111111111110000000000000000;
7'd038:bitmap<=160'b1111111111111111111111111111111111111011110000011111111111111111011111111111111111111111111111111111111111111111111111111100111111111111111111000000010000000000;
7'd039:bitmap<=160'b1111111111111111111111111111111111111111110000111111111111111111110111111111111111111111111111111111111111111111111111111001111111111111111110000100100000000000;
7'd040:bitmap<=160'b1111111111111111111111111111111111110111100110111111111111111111111101111111111111111111111111111111111111111111111111110011111111111111110000000000000000000000;
7'd041:bitmap<=160'b1111111111111111111111111111111111110111100011111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111010000000000000000000000;
7'd042:bitmap<=160'b1111111111111111111111111111111111101111100111111111111111111111111111100000111111111111111111111111111111111111111111111111111111111111110111100000000000010000;
7'd043:bitmap<=160'b1111111111111111111111111111111000001111000111111111111111111111001111100000011111111111111111111111111111111111111111111111111111111111100010001100000000011000;
7'd044:bitmap<=160'b1111111111111111111111111110111111011111000111111111111111111111111111000000000111111111111111111111111111111111111111100111111111111111000000000011000000000000;
7'd045:bitmap<=160'b1111111111111111111111111111111110111110001111111111111111111111111110000000000111111111111111111111111111111111111101101111111111111110000000000000100000010000;
7'd046:bitmap<=160'b1111111111111111111111111111111110111110001111111111111111111111111110000000000011111111111111111111111111111111111111011111111111111000000000000000010000000000;
7'd047:bitmap<=160'b1110011111111111111111011111111101111110001111111111111111111111111100000000000011111111111111111111111111111111111000011111111110000000000000000000000110000000;
7'd048:bitmap<=160'b1111001111111111111111000011111101111101001111111111111111111111111000000000000011111111111111111111111111111111100000111111111111010000000000000000000000000000;
7'd049:bitmap<=160'b1001001111111110000111000000111011111101100111111111111111111111111000000000000011111111111111111111111111111111000001111111111110000000000000000000000000001000;
7'd050:bitmap<=160'b0100101111111100000000111001111111111101001111111111111111111110010000000000000001111111111100011111111111111111001101111111110110000000000000000000000000000011;
7'd051:bitmap<=160'b0101001000000100000011111011110111110011001111111111111111111100000000000000000000111111110000001110111111111110011111111111000000000000000000000000000000010100;
7'd052:bitmap<=160'b0000000101000000000001000011110111110010001111111111111111111100000000000000000000000110101100001011111111111110001100111100000000000000000000000000001101001000;
7'd053:bitmap<=160'b0100000000000000000001100000101111110110001111111111111110111000000000000000000000000000000111000111111111111110001100111000000000000000000000000000000000000000;
7'd054:bitmap<=160'b0000000000000001000001000010001101110000001111111111111110111100000000000000000000000000001111100011111111111100000000010000000000000000000000000000000000000000;
7'd055:bitmap<=160'b0010000000000000000000000100000011110000000000001111111111000100000000000000000000000000001111100001111111111001111111100110000000000000000000000000000000000000;
7'd056:bitmap<=160'b0000000000001000000010000000000000110000000000000111111110001000000000000000000000000000001111100000111111110111111111111111000000000000000000000000000000000000;
7'd057:bitmap<=160'b0000000000000000000000000000010000000000000000000011111111100100000000000000000000000000011111110010111110001111111111001110000000000000000000000000000000000000;
7'd058:bitmap<=160'b0000000000000000100000000100000100000000000000000011111111100000000000000000000000000000000010111110011100011111111111111101000000000000000000000000000000001000;
7'd059:bitmap<=160'b0000000000000000000000000000000000000100000000000111111100000000000000000000000000000000000000011111000000011110111111111001100000000000000000000000000000000000;
7'd060:bitmap<=160'b0000000000000000000000101011000000000000000000001111111110000000000000000001100000000000000000011110100100011000011111111000100000000000000000000000000000000000;
7'd061:bitmap<=160'b0000010100000000111111111111000000100000000000000111111111100000000000000001100000000000000000011001000000010000001110110000100000000000000000000000000000000000;
7'd062:bitmap<=160'b0000000000000001011011111111000011100100111110001111111111110000000000000011100000000000000000000000000000110000011011110111110000000000000000000000000000000000;
7'd063:bitmap<=160'b0000000000000001011111111100000000001001111111001111111111110000000000000001100000000000000000000000000000111000011111110011110000000000000000000000000000000000;
7'd064:bitmap<=160'b0000000000001000111111111100000000000000111111110111111111100000000000010011100000000001000000000000000000110000011001100000110000000000000000000000000000000000;
7'd065:bitmap<=160'b0000000000011100001111111000000000000000001110000111111110100000000000010000000000000000000000000000000000010000011001100000110000100000000000000000000000000000;
7'd066:bitmap<=160'b0000000000011111011111111000000000000001000100010111111100000000000000111011000000000000000000010011110000011000011001100001100000000000000000000000000000000000;
7'd067:bitmap<=160'b0000000000111111111111111000000000000001000110100111111100000000000000001110000000000001000000000111111000011000011001100000100000000000000000000000000000000000;
7'd068:bitmap<=160'b0000000001101111111111110000000000000000000000000011111111100000000000011100000000000011000000000111111110111000011001000000101000000000000000000000000000000000;
7'd069:bitmap<=160'b0000000000111111111111100000000000000000000000000000111111110011100000011100001110000011000110000001111100001000001001000000100000000000000000000000000000000000;
7'd070:bitmap<=160'b0000010011111111111111100000011111111000000000000001111111111111010000001100011110000111100101000001001100001000001000000000100000000000000000000000000000000000;
7'd071:bitmap<=160'b0000000111111111111111000111111111111111000000000001111111111101000000001110111100000011100000000000110000001000011001000000100000000000000000000000011000000000;
7'd072:bitmap<=160'b0000011111111111111110001111111111111111110000000001111111111100000000000111111100000000100000000000110000011000011001100000110000000000000000000000011000000000;
7'd073:bitmap<=160'b0001111111111111110000011111111111111111111000000011111111110000000000000111111110000011100000000000000000011000011111100000110000000000000000000000000000000000;
7'd074:bitmap<=160'b0111111111111111000000111111111111111111111110000011111111111111000000000111111111000001100000001000000000011100111111100000111000000000000000000011000000000000;
7'd075:bitmap<=160'b0000000000000000000001111111111111111111111001100001101111111110000000000011111111100000000000000100000000011000011010100000110000000000000000000111111000000000;
7'd076:bitmap<=160'b0000000000000000000011111111111111111111110000000000000000000000000101000000111111000001000000001000000000001011111111101100110000000000000100000111110000000000;
7'd077:bitmap<=160'b0000000000000000000111111111111111111111000000000111000000000000000000000000000000000001110000000001100000001111111111111111111000000000000110011111110100000000;
7'd078:bitmap<=160'b0000000000000000000011011111111111111000000000000000000000000000000000000000000000000010010000001011100000001111111100111111111110000000000000111111100000000011;
7'd079:bitmap<=160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000010010000011000000000000110000001000000011111100000000000011111000000000011;
7'd080:bitmap<=160'b0000000000000000000000000000000000000000000000000000001110110000000000000000000000000010010000011110001000000100000011100000000110111111111111011110000000000001;
7'd081:bitmap<=160'b0000000000000000000000000000000000000000000000000000001110000000000000000000000000000110001000011111101110100000000000000000000001100010000101111000000000000000;
7'd082:bitmap<=160'b0000000000000000000000000000000000000000000000000000001110000000000000100000000000000001110000010011100110110100000001100000000000000000000011001000110000000000;
7'd083:bitmap<=160'b0011000000000000000000000000000000000000000000000000001110100000000000000000000001000000000000110110000111011111111000000000001110001001011011100100000000000000;
7'd084:bitmap<=160'b1111000000000000000000000000000000000000000000000000001100000001000000000001101000000010000000000000000000001000000000110000000000000000100000100100000000000000;
7'd085:bitmap<=160'b1111111100000000000000000000000000000000000000000000011111110000000000000011111000000010000000000000000100000000000100100000001000001000000001101011000000000000;
7'd086:bitmap<=160'b0100110100000000000000000000000000000000000000000001111111111111100000001111110000000000000000000000000000000000000000000000000000110110000011010100000000000000;
7'd087:bitmap<=160'b0000010000000000000000000000000000000000000000000001001111111100000000111111100000000000000000010000000000000000000001000000000000100000000000101000000000000000;
7'd088:bitmap<=160'b0000001000000000000000000000000000000000000000001111111111111000000111111011100000000000001000000000000000000000000011111010000000011000000000011000000000000000;
7'd089:bitmap<=160'b0000000000000000000000000000000000000000000000001111111111111011110111111000000000000000000000000000000000000000001111000001000011111000000000000000000000000000;
7'd090:bitmap<=160'b0000000000000000000000000000000000000000000000001111111111111100000000011101000000000000000011110000000000000000000110000011100010000000000100100000000000000000;
7'd091:bitmap<=160'b0000000000000000000000000000000000000000000000111111111111111111111100111111000000000000000111110000000000000000001000000011100000110000000000000000000000000000;
7'd092:bitmap<=160'b0000000000000000000000000000000000000000000011000111111111111111111001111110000000000000001100100000000000000000000000000000010000000000000101101000000000000000;
7'd093:bitmap<=160'b0000000000000000000000000000000000001100000000001111111111111111111111111111000000000111110000100000000000000000000100111100000000000000000001110000000000000000;
7'd094:bitmap<=160'b0000000000000000000000000000000000000000000000000111111111111111111111111111100000000000110010011101000000000000000001100000000000000000000000000100110000000000;
7'd095:bitmap<=160'b0000000000000000000000000000000000000000000000001011111111111111111111111111110000101000011111001010000000000000000111100111000000000000000000001000010100000000;
7'd096:bitmap<=160'b0000000000000000000000000000000000000000000000000111111111111111111111111111111000000000001111000110000000000000000000000000000000000000000000010000001000000000;
7'd097:bitmap<=160'b0000000000000000000000000000000000000000000000000111111111111111111111111111001000000000001111111101000000000000000000000000000000000000000000000000001110000000;
7'd098:bitmap<=160'b0000000000000000100000000000000000000000000000000011111111111111111111111011110000000000000000110001000000000000000000000000000000000000000000000000000011100000;
7'd099:bitmap<=160'b0000000000000000000000000000000000000000000000000111111111111111111111110100100110000000001011111000000000000000000000000000000000000000000000000000000001100000;
7'd100:bitmap<=160'b0000000000000000000000000000000000000000000000000101111111111111111111111111111100000000001101110000000000000000000000010001100000000000000000000000000000000000;
7'd101:bitmap<=160'b0000000000000000000000000000000000000000000000000001111111111111111111111111111000000000001001100000000000000000000000010000010000000000000000000000100000000000;
7'd102:bitmap<=160'b0000000000000000001111000000000000000000000000000001111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd103:bitmap<=160'b0000000000000000001110000000000000000000000000010011111111111111111111111111111100110000000000000000000000000000000010000000000000000000100001000000000000000000;
7'd104:bitmap<=160'b0000000000000000000100000000000000001000000000000000111010111111111111111111111111111111100000000100000000000000000010000000100010010000000000000000000000000000;
7'd105:bitmap<=160'b0000000000000000000000000000000000000000000000001000001111111111111111111111111111111111111101000000001000010000111111000000000000100000000000000000000000000000;
7'd106:bitmap<=160'b0000000000000000000000000000000000000000000000100000101111111111111111111111111111111111111111111110000001000001111111111000000011000000000000000000000000000000;
7'd107:bitmap<=160'b0000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111100111111111111111110000010000000000000000011100000010011;
7'd108:bitmap<=160'b0000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111010110000000000000011000011111111;
7'd109:bitmap<=160'b0000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010000000011111111111111;
7'd110:bitmap<=160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd111:bitmap<=160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd112:bitmap<=160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd113:bitmap<=160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd114:bitmap<=160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd115:bitmap<=160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd116:bitmap<=160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd117:bitmap<=160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd118:bitmap<=160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd119:bitmap<=160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
		
		endcase
	end
endmodule

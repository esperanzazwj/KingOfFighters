`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:15:54 01/08/2016 
// Design Name: 
// Module Name:    bg_rom_r 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module bg_rom_r(input wire clk, input wire[6:0] addr, output reg[159:0] bitmap);
	reg [6:0] addr_reg;
	always @(posedge clk)
		addr_reg<=addr;
	always @(*)
	begin
		case (addr_reg)
7'd000:bitmap<=160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000;
7'd001:bitmap<=160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000;
7'd002:bitmap<=160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011000;
7'd003:bitmap<=160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000;
7'd004:bitmap<=160'b0000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000;
7'd005:bitmap<=160'b0000000000000000000000000000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000;
7'd006:bitmap<=160'b0000000001000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111;
7'd007:bitmap<=160'b0000000011100000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111;
7'd008:bitmap<=160'b0000000000000000000000000000000000000000001111101111101100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110;
7'd009:bitmap<=160'b0000000000000000000000000000000000000000001111111111101110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110;
7'd010:bitmap<=160'b0000000000000001010000000000000000000000000101101101010111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111110;
7'd011:bitmap<=160'b0000000000000000000100000000000000000000000101000000110111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111101111111111111;
7'd012:bitmap<=160'b0000000000000001011110000000000000000000001100000000010110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111;
7'd013:bitmap<=160'b0000000000000000011111100000000000000000000010000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000111111101111001010000;
7'd014:bitmap<=160'b0000000000000000000111111000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111110111110100000000;
7'd015:bitmap<=160'b0000000000000000001101111110000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111010000000000000;
7'd016:bitmap<=160'b0000000000000000000001110111000000000000000011000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111000000000000000001;
7'd017:bitmap<=160'b0000000000000000000001111111110000000000000111000011111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111;
7'd018:bitmap<=160'b0000000000000000000000001110111000000000000000000011110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111;
7'd019:bitmap<=160'b0000000000000000000000000111111110000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111011;
7'd020:bitmap<=160'b0000000000000000000000000001111111100000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111;
7'd021:bitmap<=160'b0000000000000000000000000000011111110000000100000111000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111;
7'd022:bitmap<=160'b0000000000000000000000000000000111111000001110001111000000000000000010000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111;
7'd023:bitmap<=160'b0000000000000000000000000000000001111110000011001110000000000000001111000000000000000000000000000000000000000000000000000000000000000111111111100011111111111111;
7'd024:bitmap<=160'b0000000000000000000000000000000000011111100000011110000000000000111111100111000000000000000000000000000000000000000000000000000000010000000000000111111111111111;
7'd025:bitmap<=160'b0000000000000000000000000000000000000111110000011100000000000001111111111111100000000000000000000000000000000000000000000000000000000000000000000111111111111111;
7'd026:bitmap<=160'b0000000000000000001100000000000000000001100010001000000000000001111111111111100000000000000000000000000000000000000000000000000000000000000000011111111111111111;
7'd027:bitmap<=160'b0000000000000001111111100000000000000000001111010000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000111111111111111111;
7'd028:bitmap<=160'b0000000001000111111111111110000000000001000000100000000000000001111011111111111000000000000000000000000000000000000000000000000000000000000001111111111111111111;
7'd029:bitmap<=160'b0000011111111111111111111100000000000000010000100000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000001111111111111111111;
7'd030:bitmap<=160'b0000001111111111111000000000000000000000010000010000000000000000000111111111110000000000000000000000000000000000000000000000000000000000000001111111011111111110;
7'd031:bitmap<=160'b0000000000000000000000000000000000000000010010000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000001111110010111111011;
7'd032:bitmap<=160'b0000000000000000000000000000000000000000110100000011000000000000000000000000000000000000000000000000000000000000000000000000000000000000110111111111000000110111;
7'd033:bitmap<=160'b0000000000000000000000000000000000000000011000000111110100000000000000000000000000000000000000000000000000000000000000000000000111000000000011111111001000011111;
7'd034:bitmap<=160'b0000000000000000000000000000000000000000011100000011111100000000000000000000000000000000000000000000000000000000000000000000011000000000000000110110000000010101;
7'd035:bitmap<=160'b0000000000000000000000000000111111000000111000001100111111000000000000000000000000000000000000000000000000000000000000000000101000000000100000110100000000000011;
7'd036:bitmap<=160'b1111111000000000000000000011111111100001111000000001011111110000000000000000000000000000000000001100000001111111000000000010000000000001100001110000000000000000;
7'd037:bitmap<=160'b1111111100000000000000001111111111110101111100000000000111111100000000000000000000000000000000011110000011111111000000000011000000000011111011010000000000000000;
7'd038:bitmap<=160'b1111111111111000000011111111111111111011110000000000000001111111000000000000000000000000000000111111000011111111000000000000000000001011111101000000010000000000;
7'd039:bitmap<=160'b1111111111111110000111111111111111111111111100000000000000111111110000000000000000000000000111111111000111111111100000000000000000000100011110000100000000000000;
7'd040:bitmap<=160'b0111111111111101111111111111111111110111100110000000000000000111110100100000000000000000001111111111111111111111100000010000000000111000010010000000000000000000;
7'd041:bitmap<=160'b0111111111111101111111111111111111111111110000000000000000000011110110000000000000000001111111111111111111111111100001111000000011111100000000000000000000000000;
7'd042:bitmap<=160'b1000011001111111111111111111111001101111110000000000000000000000111110010000100000000001111111111111111111111111000001000011111111111001011111100000000000010000;
7'd043:bitmap<=160'b1110000000001111111111100110000000011111000011100000000000000000001100101000010000000001111111111111111111111110000111000001111111111111110111111100000000011000;
7'd044:bitmap<=160'b1111101000000111111001111000001001011011000011100000000000000000100001110000001111011111111111111111111111111110001110000011111111111111000000111111000000000000;
7'd045:bitmap<=160'b1111111100000111111011110001111110111111000011100000000000000000000000000000010111111111111111111111001111111110010000000111111111111110000000111111100000010000;
7'd046:bitmap<=160'b1111111111111111111111111111111110111111100111111100000000000000000110000000011111111111111111111110011111111111011000001111111111011000000001110011011000000000;
7'd047:bitmap<=160'b1111111111111110111111111111111101111110000111111000000000000001000110000001001111001111111111111110011111111111111000011111111110001000000100000011111110000000;
7'd048:bitmap<=160'b1011011111111111111111000111111101101101000111111100001000000010110000000000000111000000111111111100111111111001000000011111111000011000000110011111001111110000;
7'd049:bitmap<=160'b0001001111111111100111000000111011111101000111111100000000000011010000000000000110000000001100111100111111111111000000111111110000000000000000010011111111111000;
7'd050:bitmap<=160'b0100101111111110001000011001110010111111000111111110000001000000011000000010000011100000010000011001011111111110001100111111100000000000000000000001101111110111;
7'd051:bitmap<=160'b1101001111001110000011111011110111000010000111111111000001111000010000100000000100111110010000000110111111111110111111111110000000000000000000000000000111111111;
7'd052:bitmap<=160'b1010000101111000001011000011100111111010001111111111000110100111000000000000000000010100101000001011111111111110011100111100000000000000000000000000001111101111;
7'd053:bitmap<=160'b0100000010000100000001100001101011100110001111111111111110111000000000000000000000000000000110000100111111111110001110011000000000000000001000000000000000000000;
7'd054:bitmap<=160'b0110000000000001100001000011011100010100001111111111111100111100000000000000000000011000000111000000011111111000000000000001100000000000000000000000000000000000;
7'd055:bitmap<=160'b0110000000000011000000000100000011000100010000111111111100000100000000000000000010000000001011000000111111111000111111101111110000000000000110000000000000000001;
7'd056:bitmap<=160'b0000000000001001100110000000101000110000000000111111110000001000000000000000000000000010001111000000011110100111111111111111010000000000000000000000000000000010;
7'd057:bitmap<=160'b1000000000001001000010000000010011100000000000000010101011101100000000000000000000000000000110110000011110001111111111101110100000000000001100000000000000000100;
7'd058:bitmap<=160'b0000000000001100100000000100001110110010000000000001100101000000000000000000000000000000000000011000001000001001111110111101000000000000000000000000000000001000;
7'd059:bitmap<=160'b1000010000000010000000000000010010000100001110000100101000000000000000000000000000000000000000001111000000001100111111111001100000000000000000000000000000000000;
7'd060:bitmap<=160'b0000001000100100000000101000000000010001000011001000010100000000000000000001100000000000000000000000100000011000011110111000100000000000000000000000000001000000;
7'd061:bitmap<=160'b0000010100100000111001000000000000000000000100000100010100000000000000000011100000000000000000000000000000010000001000111000000000000000000000000000000100000000;
7'd062:bitmap<=160'b0000001001000000000000000000000000000100111110001000001001000000000000000011100000000000000000000000000000010000011011110111110000000000000000000000000100000000;
7'd063:bitmap<=160'b0000001110000000000000000000000000001001111111001010000010000000000000010001100000000000000000000000000000110000011001110011110000000000000000000000000000000000;
7'd064:bitmap<=160'b0000000010000000000000000000000000000001111111110000110000000000000000000011100000000000000000000000000000110000001001100000110000000000000000000000010000000000;
7'd065:bitmap<=160'b0000000000001000000000010000001000000000011111000000000000000000000000000000000000000000000000000000000000010000011000100000100000000000000000000000000000000000;
7'd066:bitmap<=160'b0000000000000000000000000000110110000011101110111000000000000000000000000011000000000000000000010000000000010000011001000000100000000000000000000000000000000000;
7'd067:bitmap<=160'b0000000000000000000000000000100000000111111111111000000000000000000000000010000000000000000000000000000000011000011001000000000000000000000000000000000000000000;
7'd068:bitmap<=160'b0000000001000000000000000000000000000000000010010011100001000000000000000000000000000000000000000000001010111000001001000000100000000000000000000000000000000000;
7'd069:bitmap<=160'b0000000000000000000000000000000000000000000100000000000000000001000000000000000000000001000000000000000010000000000000000000000000000000000000000000000000000000;
7'd070:bitmap<=160'b0000000000000000010000000000001010110000000000000000010001000101010000000000000000000111100000000001000000000000000000000000000000000000000000000000000000000000;
7'd071:bitmap<=160'b0000000001101101000000000000111100011100000000000001000111000101110000000000000000000000100000000000110000001000001000000000000000000000000000000000011000000000;
7'd072:bitmap<=160'b0000000000000000000000000000000001000110000000001000010001100110000000000000000000000000100000000000110000011000001001000000100000000000000000000000011000000000;
7'd073:bitmap<=160'b0000000000000000000000000010000000000000000000001000000000000000000000000000000000000011100000000000000001011000011111100000110000000000000000000000000000000000;
7'd074:bitmap<=160'b0000000000000000000000000000000001000010000100001000110001100001000000000000000000000011100000001000000001111000011111100000111000000000000000000011000000000000;
7'd075:bitmap<=160'b0000000000000000000000000000000100000000000000001110100000001000000000000000000001000000000000000100100001111000000010100000110000000000000000000111111000000000;
7'd076:bitmap<=160'b0000000000000000000000000000000000110000000000001000010000000000000101000000000000000011000000001100100000001011110101100100110000000000000100000111111000000000;
7'd077:bitmap<=160'b0000000000000000000000000000000000000000000000000000001111000000000000000000000000000001110000000001100000001111111111111111111000000000000110011111111100000000;
7'd078:bitmap<=160'b0000000000000000000000000000000000000000000000000000001111000000001101000000000000000010010000001011100000001111111100111111111110000000000001111111111100000000;
7'd079:bitmap<=160'b0000000000000000000000000000000000000000000000000000000000000000000110100000000000000010010000011001000000000111111011111111111111100000000011011111111000000000;
7'd080:bitmap<=160'b0000000000000000000000000000000000000000000000000000011110110000011111110000000000000010010000011111101000001111111111101111111111111111111111111111110000000000;
7'd081:bitmap<=160'b0000000000000000000000000000000000000000000000000000001110100000000000000000000000001111101000011111101110100100100011100000111111100011101111110011100000000000;
7'd082:bitmap<=160'b0000000000000000000000000000000000000000000000000000001110100000001111101000000000000111110000011111100111110110011011110011000100110000000011111000110000000000;
7'd083:bitmap<=160'b1111000000000000000000000000000000000000000000000000011110100000000000000000000000000011000000111111001111111111111111111111111111101111111111111100000000000000;
7'd084:bitmap<=160'b1111100000000000000000000000000000000000000000000100001110001001000000000001100000000000000000000000000000111110111110111100001111011111111111111100000000000000;
7'd085:bitmap<=160'b1111111100000000000000000000000000000000000000000110011111111111000001000011111000000000000000000000000100000000111111111111111111101111011111111110000000000000;
7'd086:bitmap<=160'b1111111100000000000000000000000000000000000000001101010111111111100000011111110000000000000000000000000000000011111111111100111111111111001111111110000000000000;
7'd087:bitmap<=160'b1111111010000000000000000000000000000000000000001100001111111100000000111111100000000000000000000000000000000000011111110100011111110000000101111010000000000000;
7'd088:bitmap<=160'b0000111000000000000000000000000000000010000010001111111111111010111111111111100000000000000000000000000000000000001111111011100110111000000011111100000000000000;
7'd089:bitmap<=160'b0000110000000000000000000000000000000010000010001111111111111011111110001111100000000000000000000000000000000000001111100011100011111000000011110000000000000000;
7'd090:bitmap<=160'b0000000000000000000000000000000000000110010010011111111111111111000000011111000000000000000001100000000000000000000110000011110010000000000110110000000000000000;
7'd091:bitmap<=160'b0000000000000000000000000000000000000110011110111111111111111111111100011111000000000000000001110000000000000000000000000011111000000000000000000000000000000000;
7'd092:bitmap<=160'b0000000000000000000000000000000000000011111111111111111111111111111001111110000000000000000000100000000000000000000000000000010000000000000101101000000000000000;
7'd093:bitmap<=160'b0000000000000000000000000000000011111111111111111111111111111111111111111111000000000000100000100000000000000000000000011100000000000000000000110000000000000000;
7'd094:bitmap<=160'b0000000000000000000000000000000011011111111111111111111111111111111111111111100000000000110000011100000000000000000000100000000000000000000000000100010000000000;
7'd095:bitmap<=160'b0000000000000000000000000010100011001111111110001001111111111111111111111111110000100000011110001010000000000000000111110111000000000000000000001000000000000000;
7'd096:bitmap<=160'b0000000000000000011000000100100011000000000000001111111111111111111111111111011000000000001111000110000000000000000000000000000000000000000000010000011000000000;
7'd097:bitmap<=160'b0000000000000000111100000000000011000000000000001111111111111111111111111100001000000000001111111100000100000000000000000001000000000000000000000000001110000000;
7'd098:bitmap<=160'b0000000000000000101100000000000011000000000000001111111111111111111111111000000000000000000001110000000000000000000000000000000000000000000000000000000111100000;
7'd099:bitmap<=160'b0000000000000000001000000000000011000000000000001111111111111111111111110000000110000000001111111000000000000000000000000000000000000000000000000000000000100000;
7'd100:bitmap<=160'b0000000000000000000001100000000011000000000000001101111111111111111111111111111100000000001111110000000000000000000000110011100000000000000000000000000000000000;
7'd101:bitmap<=160'b0000000000000000000010110000000011000000000000000001111111111111111111111111111000000000000001100000000000000000000000010011010000000000000000000000100000000000;
7'd102:bitmap<=160'b0000000000000000001111111000000001100000000000000001111111111111111111111111111100000000000000000000000000000000000000100101110000000000000000000000000000000010;
7'd103:bitmap<=160'b0000000000000000011111111100000001100100100000010001111111111111111111111111111100111100000100000000000000000000000111110111111011100000100001000000000000011101;
7'd104:bitmap<=160'b0000000000000000001100000100000000001100100001000000111111111111111111111111111111111111100000000111000000000101111111111111110111110000000000000001011111111011;
7'd105:bitmap<=160'b0000000000000000000011000111000000000000100000001001111111111111111111111111111111111111111111100000011101010111111111111000000111111000000000010001111111111111;
7'd106:bitmap<=160'b0000000000000000000100000111100000000000100000111101111111111111111111111111111111111111111111111111111111111111111111111111100011001111111111111111100111111111;
7'd107:bitmap<=160'b0000000000000000000000000111110001000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111111111111111111111111;
7'd108:bitmap<=160'b0000000000000000000000001111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd109:bitmap<=160'b0000000000000000000000000111111000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
7'd110:bitmap<=160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd111:bitmap<=160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd112:bitmap<=160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd113:bitmap<=160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd114:bitmap<=160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd115:bitmap<=160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd116:bitmap<=160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd117:bitmap<=160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd118:bitmap<=160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
7'd119:bitmap<=160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

		endcase
	end
endmodule
`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    21:08:34 12/11/2015 
// Design Name: 
// Module Name:    FSM_Control 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module FSM_Control(input wire clk, input wire btn, input wire[3:0] hit, 
	input wire over, input wire timeout, output wire[15:0] blood_dec, output wire ifbegin, 
	output wire reset, output wire[1:0] graph_state);
	

endmodule

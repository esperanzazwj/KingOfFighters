`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:20:47 01/05/2016 
// Design Name: 
// Module Name:    p1_rom_blue 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module p1_rom_blue(input wire clk, input wire[9:0] addr, output reg[15:0] bitmap);
//������ͼROM��16*16
reg [9:0] addr_reg;
	always @(posedge clk)
		addr_reg<=addr;
	always @(*)
	begin
		case (addr_reg)
//stay_blue&green0
10'o0000:bitmap<=16'b1111110000111111;
10'o0100:bitmap<=16'b1111100000011111;
10'o0200:bitmap<=16'b1111110000111111;
10'o0300:bitmap<=16'b1111000000011111;
10'o0400:bitmap<=16'b1100000000011100;
10'o0500:bitmap<=16'b0001100000010001;
10'o0600:bitmap<=16'b1000110000000111;
10'o0700:bitmap<=16'b1111100000011111;
10'o1000:bitmap<=16'b1111100000111111;
10'o1100:bitmap<=16'b1111000000011111;
10'o1200:bitmap<=16'b1111000000001111;
10'o1300:bitmap<=16'b1110000110000111;
10'o1400:bitmap<=16'b1110001111000011;
10'o1500:bitmap<=16'b1100011111100011;
10'o1600:bitmap<=16'b0000111111100001;
10'o1700:bitmap<=16'b0000111111110000;
//stay_blue&green1
10'o0001:bitmap<=16'b1111110000111111;
10'o0101:bitmap<=16'b1111100000011111;
10'o0201:bitmap<=16'b1111110000111111;
10'o0301:bitmap<=16'b1111000000011111;
10'o0401:bitmap<=16'b1100000000011100;
10'o0501:bitmap<=16'b0001100000010001;
10'o0601:bitmap<=16'b1000110000000111;
10'o0701:bitmap<=16'b1111100000011111;
10'o1001:bitmap<=16'b1111100000111111;
10'o1101:bitmap<=16'b1111000000011111;
10'o1201:bitmap<=16'b1111000000001111;
10'o1301:bitmap<=16'b1110000110000111;
10'o1401:bitmap<=16'b1110001111000011;
10'o1501:bitmap<=16'b1100011111100011;
10'o1601:bitmap<=16'b0000111111100001;
10'o1701:bitmap<=16'b0000111111110000;
//stay_blue&green2
10'o0002:bitmap<=16'b1111110000111111;
10'o0102:bitmap<=16'b1111100000011111;
10'o0202:bitmap<=16'b1111110000111111;
10'o0302:bitmap<=16'b1111000000011111;
10'o0402:bitmap<=16'b1100000000011100;
10'o0502:bitmap<=16'b0001100000010001;
10'o0602:bitmap<=16'b1000110000000111;
10'o0702:bitmap<=16'b1111100000011111;
10'o1002:bitmap<=16'b1111100000111111;
10'o1102:bitmap<=16'b1111000000011111;
10'o1202:bitmap<=16'b1111000000001111;
10'o1302:bitmap<=16'b1110000110000111;
10'o1402:bitmap<=16'b1110001111000011;
10'o1502:bitmap<=16'b1100011111100011;
10'o1602:bitmap<=16'b0000111111100001;
10'o1702:bitmap<=16'b0000111111110000;
//stay_blue&green3
10'o0003:bitmap<=16'b1111110000111111;
10'o0103:bitmap<=16'b1111100000011111;
10'o0203:bitmap<=16'b1111110000111111;
10'o0303:bitmap<=16'b1111000000011111;
10'o0403:bitmap<=16'b1100000000011100;
10'o0503:bitmap<=16'b0001100000010001;
10'o0603:bitmap<=16'b1000110000000111;
10'o0703:bitmap<=16'b1111100000011111;
10'o1003:bitmap<=16'b1111100000111111;
10'o1103:bitmap<=16'b1111000000011111;
10'o1203:bitmap<=16'b1111000000001111;
10'o1303:bitmap<=16'b1110000110000111;
10'o1403:bitmap<=16'b1110001111000011;
10'o1503:bitmap<=16'b1100011111100011;
10'o1603:bitmap<=16'b0000111111100001;
10'o1703:bitmap<=16'b0000111111110000;
//forward_cross_g&b0
10'o0010:bitmap<=16'b1111110000111111;
10'o0110:bitmap<=16'b1111100000011111;
10'o0210:bitmap<=16'b1111110000111111;
10'o0310:bitmap<=16'b1111110000011111;
10'o0410:bitmap<=16'b1111100000011111;
10'o0510:bitmap<=16'b1111100000011111;
10'o0610:bitmap<=16'b1111110000111111;
10'o0710:bitmap<=16'b1111100000000111;
10'o1010:bitmap<=16'b1111100000111111;
10'o1110:bitmap<=16'b1111100000001111;
10'o1210:bitmap<=16'b1111000010000111;
10'o1310:bitmap<=16'b1110000111000111;
10'o1410:bitmap<=16'b1110001111100011;
10'o1510:bitmap<=16'b1100011111000111;
10'o1610:bitmap<=16'b0000111110000111;
10'o1710:bitmap<=16'b0000111100001111;
//forward_cross_g&b1
10'o0011:bitmap<=16'b1111110000111111;
10'o0111:bitmap<=16'b1111100000011111;
10'o0211:bitmap<=16'b1111110000111111;
10'o0311:bitmap<=16'b1111110000011111;
10'o0411:bitmap<=16'b1111100000011100;
10'o0511:bitmap<=16'b1111000000011001;
10'o0611:bitmap<=16'b1100000000000111;
10'o0711:bitmap<=16'b1111000000011111;
10'o1011:bitmap<=16'b1111100000111111;
10'o1111:bitmap<=16'b1111100000111111;
10'o1211:bitmap<=16'b1111100000111111;
10'o1311:bitmap<=16'b1111100000111111;
10'o1411:bitmap<=16'b1111100000111111;
10'o1511:bitmap<=16'b1111100000111111;
10'o1611:bitmap<=16'b1111100000111111;
10'o1711:bitmap<=16'b1111100000111111;
//forward_cross_g&b2
10'o0012:bitmap<=16'b1111110000111111;
10'o0112:bitmap<=16'b1111100000011111;
10'o0212:bitmap<=16'b1111110000111111;
10'o0312:bitmap<=16'b1111110000011111;
10'o0412:bitmap<=16'b1111100000011100;
10'o0512:bitmap<=16'b1111000000011001;
10'o0612:bitmap<=16'b1100000000000111;
10'o0712:bitmap<=16'b1111000000011111;
10'o1012:bitmap<=16'b1111100000111111;
10'o1112:bitmap<=16'b1111100000111111;
10'o1212:bitmap<=16'b1111100000111111;
10'o1312:bitmap<=16'b1111100000111111;
10'o1412:bitmap<=16'b1111100000111111;
10'o1512:bitmap<=16'b1111100000111111;
10'o1612:bitmap<=16'b1111100000111111;
10'o1712:bitmap<=16'b1111100000111111;
//forward_cross_g&b3
10'o0013:bitmap<=16'b1111110000111111;
10'o0113:bitmap<=16'b1111100000011111;
10'o0213:bitmap<=16'b1111110000111111;
10'o0313:bitmap<=16'b1111110000011111;
10'o0413:bitmap<=16'b1111100000011111;
10'o0513:bitmap<=16'b1111100000011111;
10'o0613:bitmap<=16'b1111110000111111;
10'o0713:bitmap<=16'b1111100000000111;
10'o1013:bitmap<=16'b1111100000111111;
10'o1113:bitmap<=16'b1111100000001111;
10'o1213:bitmap<=16'b1111000010000111;
10'o1313:bitmap<=16'b1110000111000111;
10'o1413:bitmap<=16'b1110001111100011;
10'o1513:bitmap<=16'b1100011111000111;
10'o1613:bitmap<=16'b0000111110000111;
10'o1713:bitmap<=16'b0000111100001111;
//backforward_cross_g&b0
10'o0020:bitmap<=16'b111111000011111;
10'o0120:bitmap<=16'b1111100000011111;
10'o0220:bitmap<=16'b1111110000111111;
10'o0320:bitmap<=16'b1111110000011111;
10'o0420:bitmap<=16'b1111100000011111;
10'o0520:bitmap<=16'b1111100000011111;
10'o0620:bitmap<=16'b1111110000111111;
10'o0720:bitmap<=16'b1111100000000111;
10'o1020:bitmap<=16'b1111100000111111;
10'o1120:bitmap<=16'b1111100000001111;
10'o1220:bitmap<=16'b1111000010000111;
10'o1320:bitmap<=16'b1110000111000111;
10'o1420:bitmap<=16'b1110001111100011;
10'o1520:bitmap<=16'b1100011111000111;
10'o1620:bitmap<=16'b0000111110000111;
10'o1720:bitmap<=16'b0000111100001111;
//backforward_cross_g&b1
10'o0021:bitmap<=16'b1111110000111111;
10'o0121:bitmap<=16'b1111100000011111;
10'o0221:bitmap<=16'b1111110000111111;
10'o0321:bitmap<=16'b1111110000011111;
10'o0421:bitmap<=16'b1111100000011100;
10'o0521:bitmap<=16'b1111000000011001;
10'o0621:bitmap<=16'b1100000000000111;
10'o0721:bitmap<=16'b1111000000011111;
10'o1021:bitmap<=16'b1111100000111111;
10'o1121:bitmap<=16'b1111100000111111;
10'o1221:bitmap<=16'b1111100000111111;
10'o1321:bitmap<=16'b1111100000111111;
10'o1421:bitmap<=16'b1111100000111111;
10'o1521:bitmap<=16'b1111100000111111;
10'o1621:bitmap<=16'b1111100000111111;
10'o1721:bitmap<=16'b1111100000111111;
//backforward_cross_g&b2
10'o0022:bitmap<=16'b1111110000111111;
10'o0122:bitmap<=16'b1111100000011111;
10'o0222:bitmap<=16'b1111110000111111;
10'o0322:bitmap<=16'b1111110000011111;
10'o0422:bitmap<=16'b1111100000011100;
10'o0522:bitmap<=16'b1111000000011001;
10'o0622:bitmap<=16'b1100000000000111;
10'o0722:bitmap<=16'b1111000000011111;
10'o1022:bitmap<=16'b1111100000111111;
10'o1122:bitmap<=16'b1111100000111111;
10'o1222:bitmap<=16'b1111100000111111;
10'o1322:bitmap<=16'b1111100000111111;
10'o1422:bitmap<=16'b1111100000111111;
10'o1522:bitmap<=16'b1111100000111111;
10'o1622:bitmap<=16'b1111100000111111;
10'o1722:bitmap<=16'b1111100000111111;
//backforward_cross_g&b3
10'o0023:bitmap<=16'b1111110000111111;
10'o0123:bitmap<=16'b1111100000011111;
10'o0223:bitmap<=16'b1111110000111111;
10'o0323:bitmap<=16'b1111110000011111;
10'o0423:bitmap<=16'b1111100000011111;
10'o0523:bitmap<=16'b1111100000011111;
10'o0623:bitmap<=16'b1111110000111111;
10'o0723:bitmap<=16'b1111100000000111;
10'o1023:bitmap<=16'b1111100000111111;
10'o1123:bitmap<=16'b1111100000001111;
10'o1223:bitmap<=16'b1111000010000111;
10'o1323:bitmap<=16'b1110000111000111;
10'o1423:bitmap<=16'b1110001111100011;
10'o1523:bitmap<=16'b1100011111000111;
10'o1623:bitmap<=16'b0000111110000111;
10'o1723:bitmap<=16'b0000111100001111;
//punch_g&b0
10'o0030:bitmap<=16'b1111000011111111;
10'o0130:bitmap<=16'b1110000001111111;
10'o0230:bitmap<=16'b1111000011111111;
10'o0330:bitmap<=16'b1111100000111111;
10'o0430:bitmap<=16'b1111100000011111;
10'o0530:bitmap<=16'b1111100000011111;
10'o0630:bitmap<=16'b1111110000111111;
10'o0730:bitmap<=16'b1111100000000111;
10'o1030:bitmap<=16'b1111100000111111;
10'o1130:bitmap<=16'b1111100000001111;
10'o1230:bitmap<=16'b1111000010000111;
10'o1330:bitmap<=16'b1110000111000111;
10'o1430:bitmap<=16'b1110001111100011;
10'o1530:bitmap<=16'b1100011111000111;
10'o1630:bitmap<=16'b0000111110000111;
10'o1730:bitmap<=16'b0000111100001111;
//punch_g&b1
10'o0031:bitmap<=16'b1111000011111111;
10'o0131:bitmap<=16'b1110000001111111;
10'o0231:bitmap<=16'b1111000011111111;
10'o0331:bitmap<=16'b1111100000111111;
10'o0431:bitmap<=16'b1111100000011111;
10'o0531:bitmap<=16'b1111100000011111;
10'o0631:bitmap<=16'b1111110000111111;
10'o0731:bitmap<=16'b1111100000000111;
10'o1031:bitmap<=16'b1111100000111111;
10'o1131:bitmap<=16'b1111100000001111;
10'o1231:bitmap<=16'b1111000010000111;
10'o1331:bitmap<=16'b1110000111000111;
10'o1431:bitmap<=16'b1110001111100011;
10'o1531:bitmap<=16'b1100011111000111;
10'o1631:bitmap<=16'b0000111110000111;
10'o1731:bitmap<=16'b0000111100001111;
//punch_g&b2
10'o0032:bitmap<=16'b1111111110000111;
10'o0132:bitmap<=16'b1111111100000011;
10'o0232:bitmap<=16'b1111111110000111;
10'o0332:bitmap<=16'b1111111000001111;
10'o0432:bitmap<=16'b1111100000000000;
10'o0532:bitmap<=16'b1111100000111111;
10'o0632:bitmap<=16'b1111110000111111;
10'o0732:bitmap<=16'b1111100000111111;
10'o1032:bitmap<=16'b1111100000111111;
10'o1132:bitmap<=16'b1111100000001111;
10'o1232:bitmap<=16'b1111000010000111;
10'o1332:bitmap<=16'b1110000111000111;
10'o1432:bitmap<=16'b1110001111100011;
10'o1532:bitmap<=16'b1100011111000111;
10'o1632:bitmap<=16'b0000111110000111;
10'o1732:bitmap<=16'b0000111100001111;
//punch_g&b3
10'o0033:bitmap<=16'b1111111110000111;
10'o0133:bitmap<=16'b1111111100000011;
10'o0233:bitmap<=16'b1111111110000111;
10'o0333:bitmap<=16'b1111111000001111;
10'o0433:bitmap<=16'b1111100000000000;
10'o0533:bitmap<=16'b1111100000111111;
10'o0633:bitmap<=16'b1111110000111111;
10'o0733:bitmap<=16'b1111100000111111;
10'o1033:bitmap<=16'b1111100000111111;
10'o1133:bitmap<=16'b1111100000001111;
10'o1233:bitmap<=16'b1111000010000111;
10'o1333:bitmap<=16'b1110000111000111;
10'o1433:bitmap<=16'b1110001111100011;
10'o1533:bitmap<=16'b1100011111000111;
10'o1633:bitmap<=16'b0000111110000111;
10'o1733:bitmap<=16'b0000111100001111;
//kick_g&b0
10'o0040:bitmap<=16'b1111110000111111;
10'o0140:bitmap<=16'b1111100000011111;
10'o0240:bitmap<=16'b1111110000111111;
10'o0340:bitmap<=16'b1111000000011111;
10'o0440:bitmap<=16'b1100000000011100;
10'o0540:bitmap<=16'b0001100000010001;
10'o0640:bitmap<=16'b1000110000000111;
10'o0740:bitmap<=16'b1111100000011111;
10'o1040:bitmap<=16'b1111100000111111;
10'o1140:bitmap<=16'b1111100000001111;
10'o1240:bitmap<=16'b1111000010000111;
10'o1340:bitmap<=16'b1110000111000111;
10'o1440:bitmap<=16'b1110001111100011;
10'o1540:bitmap<=16'b1100011111000111;
10'o1640:bitmap<=16'b0000111110000111;
10'o1740:bitmap<=16'b0000111100001111;
//kick_g&b1
10'o0041:bitmap<=16'b1111110000111111;
10'o0141:bitmap<=16'b1111100000011111;
10'o0241:bitmap<=16'b1111110000111111;
10'o0341:bitmap<=16'b1111110000011111;
10'o0441:bitmap<=16'b1111100000011100;
10'o0541:bitmap<=16'b1111000000011001;
10'o0641:bitmap<=16'b1100000000000111;
10'o0741:bitmap<=16'b1111000000011111;
10'o1041:bitmap<=16'b1111100000111111;
10'o1141:bitmap<=16'b1111100000111111;
10'o1241:bitmap<=16'b1111100000111111;
10'o1341:bitmap<=16'b0000000000111111;
10'o1441:bitmap<=16'b1111100011111111;
10'o1541:bitmap<=16'b1111100011111111;
10'o1641:bitmap<=16'b1111100011111111;
10'o1741:bitmap<=16'b1111100011111111;
//kick_g&b2
10'o0042:bitmap<=16'b1111000011111111;
10'o0142:bitmap<=16'b1110000001111111;
10'o0242:bitmap<=16'b1111000011111111;
10'o0342:bitmap<=16'b1111100000111111;
10'o0442:bitmap<=16'b1111100000011100;
10'o0542:bitmap<=16'b1111000000011001;
10'o0642:bitmap<=16'b1100000000000111;
10'o0742:bitmap<=16'b1111000000011111;
10'o1042:bitmap<=16'b1111100000111111;
10'o1142:bitmap<=16'b1111100010001111;
10'o1242:bitmap<=16'b1111100011000111;
10'o1342:bitmap<=16'b1111100011100011;
10'o1442:bitmap<=16'b1111100011110001;
10'o1542:bitmap<=16'b1111100011111000;
10'o1642:bitmap<=16'b1111100011111100;
10'o1742:bitmap<=16'b1111100011111110;
//kick_g&b3
10'o0043:bitmap<=16'b1111110000111111;
10'o0143:bitmap<=16'b1111100000011111;
10'o0243:bitmap<=16'b1111110000111111;
10'o0343:bitmap<=16'b1111110000011111;
10'o0443:bitmap<=16'b1111100000011100;
10'o0543:bitmap<=16'b1111000000011001;
10'o0643:bitmap<=16'b1100000000000111;
10'o0743:bitmap<=16'b1111000000011111;
10'o1043:bitmap<=16'b1111100000111111;
10'o1143:bitmap<=16'b1111100000111111;
10'o1243:bitmap<=16'b1111100000111111;
10'o1343:bitmap<=16'b0000000000111111;
10'o1443:bitmap<=16'b1111100011111111;
10'o1543:bitmap<=16'b1111100011111111;
10'o1643:bitmap<=16'b1111100011111111;
10'o1743:bitmap<=16'b1111100011111111;


		
			
		endcase
	end

endmodule
